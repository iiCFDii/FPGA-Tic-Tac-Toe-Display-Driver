module shape4 (output [79:0] empty [0:79]
				  );

logic [79:0] inputImage4 [0:79] = '{   		  
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111,
80'b11111111111111111111111111111111111111111111110111111111111111111111111111111111
														  };
														  
						  
assign empty = inputImage4;
			  
endmodule
