module player2 (output [24:0] oshapes [0:24]
				  );

logic [24:0] inputImage3 [0:24] = '{   		  

25'b11111111111111111111111111,
25'b10000000000011110000000011,
25'b10111111111011111111111011,
25'b10111111111011111111111011,
25'b10111111111011111111111011,
25'b10111111111011111111111011,
25'b10111111111011111111111011,
25'b10111111111011111111111011,
25'b10111111111011111111111011,
25'b10111111111011111111111011,
25'b10000000000011111111111011,
25'b10111111111111111111111011,
25'b10111111111111110000000011,
25'b10111111111111110111111111,
25'b10111111111111110111111111,
25'b10111111111111110111111111,
25'b10111111111111110111111111,
25'b10111111111111110111111111,
25'b10111111111111110111111111,
25'b10111111111111110111111111,
25'b10111111111111110111111111,
25'b10111111111111110111111111,
25'b10111111111111110111111111,
25'b10111111111111110000000011,
25'b11111111111111111111111111
};
														  
						  
assign oshapes = inputImage3;
			  
endmodule