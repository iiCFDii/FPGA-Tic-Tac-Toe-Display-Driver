module count5 (output [24:0] oshapes [0:24]
				  );

logic [24:0] inputImage3 [0:24] = '{   		  

25'b1111111111111111111111111,
25'b1111111111111111111111111,
25'b1111111111111111111111111,
25'b1011101110111011111111111,
25'b1001101110111011111111111,
25'b1010101110111011111111111,
25'b1011001110111011111111111,
25'b1011101110111011111111111,
25'b1011100110111011111111111,
25'b1011101010111011111111111,
25'b1011101100111011111111111,
25'b1011101110111011111111111,
25'b1011101110011011111111111,
25'b1011101110101011111111111,
25'b1011101110110011111111111,
25'b1011101110111011111111111,
25'b1011101110111001111111111,
25'b1011101110111010111111111,
25'b1011101110111011111111111,
25'b1011101110111011111111111,
25'b1011101110111011111111111,
25'b1011101110111011111111111,
25'b1111111111111111111111111,
25'b1111111111111111111111111,
25'b1111111111111111111111111
};
		
														  
						  
assign oshapes = inputImage3;
			  
endmodule