module player1 (output [24:0] oshapes [0:24]
				  );

logic [24:0] inputImage3 [0:24] = '{   		  

25'b1111111111111111111111111,
25'b1000000000001111111011111,
25'b1011111111101111111011111,
25'b1011111111101111111011111,
25'b1011111111101111111011111,
25'b1011111111101111111011111,
25'b1011111111101111111011111,
25'b1011111111101111111011111,
25'b1011111111101111111011111,
25'b1011111111101111111011111,
25'b1000000000001111111011111,
25'b1011111111111111111011111,
25'b1011111111111111111011111,
25'b1011111111111111111011111,
25'b1011111111111111111011111,
25'b1011111111111111111011111,
25'b1011111111111111111011111,
25'b1011111111111111111011111,
25'b1011111111111111111011111,
25'b1011111111111111111011111,
25'b1011111111111111111011111,
25'b1011111111111111111011111,
25'b1011111111111111111011111,
25'b1011111111111111111011111,
25'b1111111111111111111111111
};
														  
						  
assign oshapes = inputImage3;
			  
endmodule