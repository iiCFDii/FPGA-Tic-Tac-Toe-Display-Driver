module shape2 (output [24:0] xshapes [0:24]
				  );

logic [24:0] inputImage2 [0:24] = '{   		  

25'b01111111111111111111111101,
25'b10111111111111111111111011,
25'b11011111111111111111110111,
25'b11101111111111111111101111,
25'b11110111111111111111011111,
25'b11111011111111111110111111,
25'b11111101111111111101111111,
25'b11111110111111111011111111,
25'b11111111011111110111111111,
25'b11111111101111101111111111,
25'b11111111110111011111111111,
25'b11111111111010111111111111,
25'b11111111111101111111111111,
25'b11111111111010111111111111,
25'b11111111110111011111111111,
25'b11111111101111101111111111,
25'b11111111011111110111111111,
25'b11111110111111111011111111,
25'b11111101111111111101111111,
25'b11111011111111111110111111,
25'b11110111111111111111011111,
25'b11101111111111111111101111,
25'b11011111111111111111110111,
25'b10111111111111111111111011,
25'b01111111111111111111111101
};
														  
						  
assign xshapes = inputImage2;
			  
endmodule