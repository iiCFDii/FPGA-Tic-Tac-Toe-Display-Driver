module shape3 (output [24:0] oshapes [0:24]
				  );

logic [24:0] inputImage3 [0:24] = '{   		  

25'b11111111000000000001111111,
25'b11111000111111111100011111,
25'b11110011111111111110011111,
25'b11110011111111111111001111,
25'b11110011111111111111001111,
25'b11110011111111111111001111,
25'b11110011111111111111001111,
25'b11110011111111111111001111,
25'b11110011111111111111001111,
25'b11110011111111111111001111,
25'b11110011111111111111001111,
25'b11110011111111111111001111,
25'b11110011111111111111001111,
25'b11110011111111111111001111,
25'b11110011111111111111001111,
25'b11110011111111111111001111,
25'b11110011111111111111001111,
25'b11110011111111111111001111,
25'b11110011111111111111001111,
25'b11110011111111111111001111,
25'b11110011111111111111001111,
25'b11110011111111111111001111,
25'b11111000111111111100011111,
25'b11111111000000000001111111,
25'b11111111111111111111111111
};
														  
						  
assign oshapes = inputImage3;
			  
endmodule