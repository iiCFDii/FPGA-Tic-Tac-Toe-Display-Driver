module count3 (output [24:0] oshapes [0:24]
				  );

logic [24:0] inputImage3 [0:24] = '{   		  

25'b1111111111111111111111111,
25'b1111111111111111111111111,
25'b1111111111111111111111111,
25'b1011101110111111111111111,
25'b1011101110111111111111111,
25'b1011101110111111111111111,
25'b1011101110111111111111111,
25'b1011101110111111111111111,
25'b1011101110111111111111111,
25'b1011101110111111111111111,
25'b1011101110111111111111111,
25'b1011101110111111111111111,
25'b1011101110111111111111111,
25'b1011101110111111111111111,
25'b1011101110111111111111111,
25'b1011101110111111111111111,
25'b1011101110111111111111111,
25'b1011101110111111111111111,
25'b1011101110111111111111111,
25'b1011101110111111111111111,
25'b1011101110111111111111111,
25'b1011101110111111111111111,
25'b1111111111111111111111111,
25'b1111111111111111111111111,
25'b1111111111111111111111111
};
		
														  
						  
assign oshapes = inputImage3;
			  
endmodule